-- Create Date:    	12:48:29 02/26/2017 
-- Design Name: 		Connect Four Display Module
-- Module Name:   	DisplayModule - Behavioral 
-- Project Name: 		Connect Four
-- Target Devices:	Nexys 4 DDR
-- Description: 		Module for the Connect Four game that implements display to a screen via VGA.
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use IEEE.STD_LOGIC_UNSIGNED.all;
use work.GamePackage.GAME_BOARD;

entity DisplayModule is
end DisplayModule;

architecture Behavioral of DisplayModule is

begin


end Behavioral;

